
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package Page_table_Type is
Type ppn_addresses is array (511 Downto 0) of std_logic_vector(6 Downto 0);
end package Page_table_Type;


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;




entity Page_table is
	port(
		virtual_address : IN std_logic_vector(15 downto 0);
		physical_address: OUT std_logic_vector(13 downto 0)
	);
end Page_table;

architecture Behavioral of Page_table is

begin
process(virtual_address, valid_bit)
	variable page_offset: std_logic_vector(6 downto 0);
	variable final_address : std_logic_vector(13 downto 0);
	variable vpn: std_logic_vector(8 downto 0);
	variable ppn: std_logic_vector(6 downto 0);
	variable my_ppn_addresses : ppn_addresses;
	variable index : Integer;
	begin
		page_offset := virtual_address(6 downto 0);
		vpn := virtual_address(15 downto 7);
		index = to_integer(unsigned(vpn));
		my_ppn_addresses := ( "1101010",    "1001011",    "1100001",    "0101010",
         "1101000",    "0010011",    "1011010",    "0010010",
         "0011001",    "0010110",    "1111101",    "0111111",
         "0010000",    "1001111",    "1110110",    "0011110",
         "1111000",    "1001000",    "0100100",    "1110101",
         "0010011",    "0100000",    "0000101",    "1011000",
         "0001110",    "0100111",    "1001110",    "0110100",
         "1010010",    "1011100",    "1111011",    "0010011",
         "0111101",    "1111101",    "0011110",    "1011001",
         "1100100",    "0110101",    "0011010",    "0011100",
         "0000010",    "1111010",    "0110011",    "0110000",
         "1001010",    "1010000",    "1010011",    "0001111",
         "1010010",    "0010001",    "1000111",    "0101011",
         "0011011",    "1010001",    "1100010",    "1101011",
         "1111001",    "0011111",    "0101100",    "0101010",
         "1000100",    "0000101",    "0111011",    "1011101",
         "1110011",    "0101100",    "0011001",    "1000010",
         "0001000",    "1100100",    "1001101",    "1110001",
         "0111101",    "0000101",    "1111010",    "1111111",
         "1111011",    "1101110",    "1011000",    "0010100",
         "0110110",    "1011110",    "0111011",    "0011100",
         "0111010",    "0001111",    "1100010",    "0010101",
         "1101110",    "1011010",    "1011000",    "1101110",
         "0011011",    "1001100",    "1101110",    "0001001",
         "0000000",    "0111111",    "0100101",    "0100001",
         "1010110",    "0110101",    "0011111",    "0011001",
         "1011101",    "0001110",    "1101110",    "1000010",
         "0100100",    "1100111",    "0000100",    "1111110",
         "1001110",    "1000011",    "0111101",    "1110011",
         "1111000",    "1100011",    "0111101",    "0111101",
         "1111110",    "1011011",    "1111110",    "0101100",
         "0110101",    "1000010",    "0000011",    "0100110",
         "0101101",    "1011010",    "1110011",    "0001101",
         "0001110",    "0010010",    "1110101",    "1000101",
         "1100101",    "0111011",    "1111110",    "0011111",
         "0100110",    "0011101",    "0100111",    "1011101",
         "1010101",    "0011011",    "0110100",    "0000110",
         "0111110",    "0110000",    "1110000",    "1000110",
         "1100100",    "1101010",    "1011101",    "1100011",
         "1110111",    "1111101",    "0010001",    "1110110",
         "1011011",    "1100001",    "1110101",    "0110111",
         "1110100",    "1111110",    "0011010",    "1110000",
         "1110100",    "0100010",    "1010000",    "0110000",
         "1010111",    "1110110",    "1111100",    "1001101",
         "1101000",    "1100101",    "1011001",    "0111010",
         "0111010",    "0111011",    "0010110",    "1011101",
         "0101001",    "0011010",    "0111001",    "0100000",
         "0011011",    "0100101",    "1000110",    "0010000",
         "0000110",    "0010101",    "1001011",    "0011110",
         "1010111",    "0000001",    "1010011",    "1010101",
         "1011100",    "1001011",    "1101011",    "1010110",
         "0010110",    "1110001",    "0000010",    "0011100",
         "1111100",    "1001001",    "0010010",    "0101111",
         "0000101",    "1110100",    "0011111",    "0010011",
         "0111010",    "1010011",    "0000110",    "0011000",
         "0110011",    "1101001",    "1111111",    "1000110",
         "1001101",    "1100000",    "1111000",    "0110001",
         "0111110",    "0100100",    "1000010",    "0001110",
         "1011001",    "0101011",    "1101110",    "1000001",
         "1000001",    "0010000",    "0010010",    "0111101",
         "0111100",    "0111100",    "1101000",    "1101100",
         "0000110",    "1100110",    "0110111",    "1010101",
         "0010101",    "0101001",    "1010001",    "1010010",
         "0001110",    "0000101",    "0001111",    "0011101",
         "1000011",    "1101000",    "1010001",    "1100011",
         "1111011",    "0100110",    "1100101",    "1000101",
         "1011001",    "1010000",    "1110110",    "0011001",
         "1101100",    "1101001",    "0011001",    "0011111",
         "0001011",    "0101011",    "1100101",    "0000101",
         "1001000",    "1100110",    "0000001",    "1101011",
         "1101111",    "0001100",    "0000010",    "0010100",
         "1101000",    "0101100",    "1001111",    "1101001",
         "0100110",    "1111101",    "0000000",    "1001010",
         "0100110",    "1111100",    "0100010",    "1011010",
         "1000100",    "1110001",    "1101011",    "1101010",
         "1001111",    "0101000",    "0111001",    "1011100",
         "0011111",    "0100111",    "1000010",    "0011110",
         "1001100",    "1000101",    "1011110",    "1011100",
         "0001011",    "0101001",    "0110110",    "1000010",
         "0111001",    "1010101",    "1000001",    "1011110",
         "0001110",    "0001101",    "1001110",    "1001010",
         "0111000",    "0101001",    "1111001",    "0010011",
         "1010101",    "1100000",    "1111110",    "1110000",
         "1100110",    "0111001",    "1110011",    "0101110",
         "0101101",    "0101010",    "1111000",    "0110100",
         "1010000",    "1111001",    "1011011",    "0100011",
         "1011111",    "0010100",    "0011011",    "0010111",
         "0111001",    "0001101",    "1011000",    "0101100",
         "1101010",    "0101110",    "0110000",    "0110100",
         "1001011",    "0101011",    "0000101",    "0111001",
         "0110100",    "0101010",    "1011000",    "0010110",
         "1101000",    "1011110",    "0011110",    "0000010",
         "0101011",    "0100010",    "1110111",    "1100101",
         "0000101",    "0100110",    "0000001",    "1100111",
         "1001010",    "1001011",    "1100001",    "1010011",
         "0111001",    "1101011",    "0111101",    "0111010",
         "1000011",    "0101101",    "0110101",    "0011110",
         "0011101",    "0000000",    "0011001",    "0110100",
         "1111111",    "1000000",    "0110111",    "1011010",
         "0110101",    "0101110",    "0010011",    "1100101",
         "0011110",    "1101000",    "1011110",    "1101101",
         "1000110",    "0101101",    "1011011",    "1011010",
         "0101100",    "1111001",    "0111010",    "0011001",
         "0110100",    "0000011",    "0100100",    "0101001",
         "1010010",    "0101101",    "1101010",    "0001001",
         "0100000",    "0011100",    "1010100",    "0000101",
         "1001011",    "0000000",    "0000111",    "1001001",
         "0001011",    "0111000",    "0000010",    "1000011",
         "0011111",    "0011101",    "1100011",    "1001110",
         "1001011",    "0001010",    "0111010",    "0010011",
         "1111101",    "1111111",    "1010111",    "1110110",
         "1001110",    "1110010",    "0101111",    "1100111",
         "1000110",    "0000101",    "1001010",    "1110000",
         "0011011",    "0110110",    "0100000",    "0101110",
         "1010110",    "0011011",    "0100111",    "1000100",
         "0011010",    "1010111",    "0111100",    "0001100",
         "1110000",    "1110010",    "0010011",    "1010100",
         "1000101",    "1010001",    "1111000",    "1011011",
         "1101101",    "1101000",    "0000010",    "0011011",
         "1010011",    "0001011",    "0100101",    "1110010",
         "1111011",    "0001111",    "0110101",    "1100101",
         "1000000",    "0100111",    "1000100",    "0010001",
         "1001100",    "0110100",    "0000011",    "1111111",
         "0001101",    "1001111",    "1011111",    "0100000",
         "0001011",    "0000111",    "0010010",    "0111101",
         "0111011",    "1000111",    "1011011",    "1001101",
         "1010101",    "1100111",    "1011000",    "1100111",
         "0000110",    "1111011",    "1111101",    "0011010");
		ppn := my_ppn_addresses(index);
		final_address(6 downto 0) := page_offset;
		final_address(13 downto 7) := ppn;
		physical_address <= final_address;
	end process
end Behavioral;





