
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.Numeric_Std.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package StorageType is
Type return_page is array (15 Downto 0) of std_logic_vector(63 Downto 0);
Type pages is array (7 Downto 0) of return_page; 
end package StorageType;




library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use work.StorageType.all;

entity Storage is
	port(
		i: IN STD_LOGIC_VECTOR(8 Downto 0);
		Output: OUT return_page);
end Storage;

architecture Behavioral of Storage is
begin
process(i)
	
	Variable input:Integer; 
	Variable Addresses: pages;
	begin 
		input := to_integer(unsigned(i));
		Addresses := 	(       
         

         ("1110111011001101011101110011000010100111000101000101111001010010",
         "0001011011101100001111111100111111110110011101100011110010001001",
         "0100100100110100010110010100101111111110110000000100001111110011",
         "1110010000001011101011010010101001010110101110010110011010001000",
         "1101010100100110100101000000100101110000110110110010010100101000",
         "1110001111011111110110110000110100101100101010010010101000011110",
         "0010011111110101100110001010000001110110010100011111100010111100",
         "0100000010100101110010110001110100111110010100110001010110100011",
         "0100011111101101011101001101011010001011010010101011101111111111",
         "0001010111011111001100010110101111011011101110101011000101011111",
         "1101101011010101110111110010001101111010000001111100110010011100",
         "1000010010101100101110010100000010000100111011001011111101001001",
         "1010000010101101001100011001111001001010101001010100100010010001",
         "1111001001110010111001110110110010111101011001111000101111101010",
         "0100001011110111101111110000000101111111101011101011100110000111",
         "1000000111011110110001111001101010110110110000111111000001111111")
			,
         ("1000111011101000000100100010110111111010000000101101110101100101",
         "1111111010101000001111000110110100111110001001100110010011110110",
         "1001101001010111000101100111111100101110010011010100111110010001",
         "0110101011000100010001101000111010001000010100001110101110000000",
         "0011110011001100110110010001010011011111011000000100001111110101",
         "0000011111111100000111110011010100101001010100111001011011000001",
         "1111110111101100110001000110100100101111011010110001100100110011",
         "0111100111010101101111101111110101010101111100101111000100110000",
         "0011100110000001111010101011100000001101010110011110011111000101",
         "0011110100111001001110110010111011100101110110101011011011111100",
         "0110011010011111001010101110101101101010100101111011101001100111",
         "0001011110101110010010101100100010101010100011000110001110001011",
         "0100101100001010100110101001000110001111000101101100010111100110",
         "1010100111111011000010010001101010110001001000111111101011000111",
         "0011110001010100111100010000000010110010101000110011011100100101",
         "1001001001011011001110111110111011110110010100001101111101001100")
			,
         ("1100110001010000110111110110000010101010010011000011110111111000",
         "0100101110111011101110111010001101011011000000001101010011110101",
         "1100001001111010100111010010001000010011010011011111100111101001",
         "1110000011000101100000111001101111101100000101111000001101110100",
         "0000010000011110001110101001110100100101001110000111001000100001",
         "0001001110011000001011001110011000100000000011010110111001001010",
         "1001000001000001100011100010101011110100111001110101100110000011",
         "0110001000010100001001000100100110111000011011101111001110111001",
         "1110100100001000100110010011111001011010011111011000001000010100",
         "0001000100000011101010101110001011001000101011011010111101100100",
         "0110001000010100111000111011011101000000110000110111010011001001",
         "1101010100110000111111001110111011100111010100001011111101111110",
         "0011001100011001011101011001110110001001111111001000000111011110",
         "1011100011011010101100001000010001001000100001110010110010100100",
         "1010111100000111001001101110100110100001011111110001011011010010",
         "0011010100111110111001101111001000000010010101101111111110110011")
			,
         ("1111100101100000010000001000111001011001010100111110101111011011",
         "0111110110100010000000011011010011111010001010011000111001100000",
         "1001110011101010010011010011100011111111000111111111011101101101",
         "0100011011010101001011001111000010101100010011110001011111100001",
         "0001111101001101001100011110001110101010100101011000111010010000",
         "0011101001100101101001011111010101101000110100011010110101111001",
         "1100100001001011110011111100010011110111010100001011100010100101",
         "0101100011000100011000010010111101110111111110000110010011101010",
         "1110001100000001111111011111001100010001101011110011111001010101",
         "1011110011111010010100000011111010111110000111011000101010111000",
         "0000010010111001001111101001111110110110001011100100001100000101",
         "1001010101101111110001010011010010000011110001101111001101010000",
         "1100010101001011001010111100011010000000010110101000011111111001",
         "1101111001110101001101100111010111110001010111111000101111011111",
         "1011111011100110010111101101010010011110001100000110011101100111",
         "1010010101010001010101001011001110100001100101010000011110001110")
			,
         ("0100110000001000010110110010101000000010111011110010001111010000",
         "0000101110101011010111011111010100100111111001001001100010000001",
         "1000000001010001011000111110001100110001111110111111010111110000",
         "1011010111110011110001000111100001000011101111101011101000001001",
         "0000000011111101111100011011011110100000001010011000011000011110",
         "0101010010100000000100011001000011001011011100101011011001110000",
         "1100010010110000101010001111011110000011010100000000100001010010",
         "0011001010001011001100000100010111111000011001010101101010000000",
         "0000100011010010000000110011010110001101010110110110001001111111",
         "1000010100011001000010111100010101111101110011111100101000000101",
         "1010100011101010101110000111011011110111011101110111010110110100",
         "1110010100010001110100000010000101101000110111011100100011011011",
         "0110100010100000110101010011111010110011011000000101001100000011",
         "1001110100000011100000111100000000000010001101110110111010001011",
         "0010010000010110111110000011011111101110011011100001101110101010",
         "1001111011100111000000011001010010000110000101000111000010110011")
			,
         ("1011111001110000101110111001000000010111101010111110000001101100",
         "0100001101000111111001010110100111110110011001100011100011110111",
         "1000100000101001100111111101100010111111000110110101011010011000",
         "1001100111111011100010000001001110100111010101010110001100011001",
         "1111110110001101101011110011011110001001011010011110100100101000",
         "0100001001010101100111000110010101111101100000101011100111111000",
         "1111011111011000001100111010110001100001010101001110111100101001",
         "1001111101001000001101011111101101101001100000101010001000111011",
         "1110110000100011001001000110110101100010000101011010101001000110",
         "1010100110010110110000100000000111011101101110011100101011010110",
         "1100011110001000110010110111101010000100000111010101100010101111",
         "1001011111011010111100100011011001101110000011101011111010100001",
         "1011100110001101110110000010001001000001010110111110100100011100",
         "1111011100011001100100111001001110110010011100110010110000011100",
         "1010010010000100101111100010111101101001101111101100110011111010",
         "0101011101110101011110111000000111101101100000000011110111000010")
			,
         ("0001110110000111001011100000010101000111101011000011101111111101",
         "0110011001100000011011000110100001100000101001100101110001110111",
         "1001001001110000001010001000000100000100111101101000110001011100",
         "0100111110000000100000101011011110110000100101001101100010111110",
         "0001110011011101010101011001011010111000010111100010011101110110",
         "0100100100101010011111110001101000101000111110010000001011111010",
         "1010000110011011100100100101011000000110011010100110101110111010",
         "0011111111100111100011000111111100100000110001110101000010101000",
         "0010111110011001010111111110001110110100100110100000110011111010",
         "1011010101101100010000101100001000000010011000000111001111010100",
         "1100010101110010001111001111010011101001000011001010101000010111",
         "0010100110010110110011000100000001001001100001110010101101000000",
         "0101000001011100000000011110000110010001000100100011111011100110",
         "1100011111101010001010001001000010110110111101010001000111111101",
         "1101110011100001100011100011101000001011111111000001110010010001",
         "1101010100110010001101010010010100110001000110111000011000110111")
			,
         ("0100100011011100011010100010110011000000110111101100101000111011",
         "1000011001111000010010101111110001100111110011001011000110010010",
         "1001101001101110011110111100001010111110111110010001110110100101",
         "1001001011101111101100001111001010110000010110001000100001010111",
         "0110000110100011001000010101001001101011001011101100100011011100",
         "0001001100110010001110010001111001000011011001010000001111100110",
         "1100000111101110111111011100101100101101100001101001111101001100",
         "0111010111010110010001101111101100010100110000111010101001001110",
         "1101011100000010101111010100110001000000100000110011011100011010",
         "1110101000010110000000000001101110110011110101010111111100011100",
         "1100010000100010010110100010000110101101100000101110100000111100",
         "0111010000011110010010010110100011000000001100111100101111110000",
         "1010100100110001100000100001110000111011000101011011000101001110",
         "0011100100101111110000011000100001101001100110101111010101010101",
         "1100110011001001010000000101001101010100011001010111101100110100",
         "1001010110110010000011110101000010001111010110111010101100100010")

			);


       
		
	
		Output <= Addresses(input);
	end process;
end Behavioral;

