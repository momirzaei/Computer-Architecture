--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   18:33:48 07/08/2022
-- Design Name:   
-- Module Name:   E:/Xilinx/Project/simulatre_processor.vhd
-- Project Name:  Project
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: Processor
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY simulatre_storage IS
END simulatre_storage;
 
ARCHITECTURE behavior OF simulatre_storage IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT storage
    PORT(
         i : IN  std_logic_vector(8 downto 0);
         Output : OUT  return_page
        );
    END COMPONENT;
    

   --Inputs
   signal i : std_logic_vector(8 downto 0) := (others => '0');

 	--Outputs
   signal Output : return_page;
   -- No clocks detected in port list. Replace <clock> below with 
   -- appropriate port name 
 
   constant clk_period : time := 10 ns;
	signal clk :std_logic;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: storage PORT MAP (
          i => i,
          Output => Output
        );

   -- Clock process definitions
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 100 ns;	
		i <= "000000000";
      wait for clk_period*10;

      -- insert stimulus here 

      wait;
   end process;

END;
